//1.Definicion del modulo y sus Ins and Outs
//Dentro del parentesis se define los I/O
module _and (input a, input b, output c);
//2.Definen cables o componentes 
//NA
//3.Asignaciones, instancias y conexiones
assign c = a & b;
endmodule